package SHARED_pkg;
    parameter FIFO_WIDTH = 16;
    parameter FIFO_DEPTH = 8 ;
    integer error_count   = 0 ;
    integer correct_count = 0 ;
    bit test_finished ;
endpackage



