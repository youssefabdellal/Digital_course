module p3 (a,b,c);
input wire [3:0] a,b ;
output wire [3:0] c ;

assign c = a + b ;
endmodule