package SHARED_pkg;
    bit test_finished;
endpackage