package shift_reg_agent_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import shift_reg_sequencer_pkg::*;
    import shift_reg_driver_pkg::*;
    import shift_reg_config_pkg::*;
    import shift_reg_monitor_pkg::*;
    import shift_reg_item_pkg::*;

    class shift_reg_agent extends uvm_agent;
        `uvm_component_utils(shift_reg_agent)
        shift_reg_sequencer sqr ;
        shift_reg_driver drv ;
        shift_reg_monitor mon;
        shift_reg_config shift_cfg;
        uvm_analysis_port #(shift_reg_item) agt_ap;

        function new(string name = "shift_reg_agent" , uvm_component parent = null );
            super.new(name, parent);
        endfunction 

        function void build_phase (uvm_phase phase);
            super.build_phase(phase);
            if (!uvm_config_db #(shift_reg_config)::get(this, "", "shift_CFG", shift_cfg)) begin
                `uvm_fatal("build_phase", "shift_reg_AGENT - unable to get configuration object");
            end 
            mon = shift_reg_monitor::type_id::create("mon",this);
            agt_ap = new("agt_ap",this);
            if (shift_cfg.is_active == UVM_ACTIVE) begin
                drv = shift_reg_driver::type_id::create("drv",this);
                sqr = shift_reg_sequencer::type_id::create("sqr",this);
            end 
        endfunction

        function void connect_phase(uvm_phase phase);
            super.connect_phase(phase);
            mon.shift_reg_vif = shift_cfg.shift_reg_vif;
            mon.mon_ap.connect(agt_ap);
            if (shift_cfg.is_active == UVM_ACTIVE) begin
                drv.seq_item_port.connect(sqr.seq_item_export);
                drv.shift_reg_vif = shift_cfg.shift_reg_vif;
            end
        endfunction
        
    endclass 
endpackage