interface shift_reg_if ();
  logic reset; 
  logic serial_in, direction, mode;
  logic [5:0] datain, dataout;
endinterface 