module shift_reg (serial_in, direction, mode, datain, dataout);
input serial_in, direction, mode;
input [5:0] datain;
output reg [5:0] dataout;

always @(*) begin
      if (mode) // rotate
         if (direction) // left
            dataout = {datain[4:0], datain[5]};
         else
            dataout = {datain[0], datain[5:1]};
      else // shift
         if (direction) // left
            dataout = {datain[4:0], serial_in};
         else
            dataout = {serial_in, datain[5:1]};
end
endmodule